# ====================================================================
#
#      hal_arm_arm9_mini2440.cdl
#
#      FriendlyARM MINI2440 evaluation board HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):	T.C. Chiu <TCChiu@sq.com.tw>
# Contributors:	T.C. Chiu <TCChiu@sq.com.tw>
# Date:		2009-12-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_ARM9_MINI2440 {
	display		"FriendlyARM MINI2440 development board"
	parent		CYGPKG_HAL_ARM_ARM9_S3C2440X
	hardware
	include_dir	cyg/hal
	define_header	hal_arm_arm9_mini2440.h
	description	"
		The MINI2440 HAL package provides the support needed to run eCos on Samsung 
		S3C2440X (ARM920T) based boards."

	compile		mini2440_misc.c

	implements	CYGINT_HAL_DEBUG_GDB_STUBS
	implements	CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
	implements	CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
	implements	CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT

	define_proc {
		puts $::cdl_header "/***** package proc output start *****/"
		puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H		<pkgconf/hal_arm.h>"
		puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H		<pkgconf/hal_arm_arm9.h>"
		puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H	<pkgconf/hal_arm_arm9_s3c2440x.h>"
		puts $::cdl_system_header "#define CYGBLD_HAL_BOARD_H		<pkgconf/hal_arm_arm9_mini2440.h>"
		puts $::cdl_header "#define CYGBLD_HAL_PLF_INTS_H		<cyg/hal/hal_platform_ints.h>"
		puts $::cdl_header "#define HAL_PLATFORM_CPU			\"ARM9\""
		puts $::cdl_header "#define HAL_PLATFORM_BOARD			\"FriendlyARM mini2440\""
		puts $::cdl_header "#define HAL_PLATFORM_EXTRA			\"\""
		puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE		1999"
		puts $::cdl_header "/***** package proc output end *****/"
	}

	cdl_component CYG_HAL_STARTUP {
		display		"Startup type"
		flavor		data
		legal_values	{ "RAM" "ROM" "ROMRAM" }
		default_value	{ "RAM" }
		no_define
		define		-file system.h CYG_HAL_STARTUP
		description	"
			When targetting the MINI2440 evaluation board it is possible to build 
			the system for either RAM bootstrap or ROM bootstrap(s). Select 
			'ram' when building programs to load into RAM using eCos GDB stubs.
			Select 'rom' when building a stand-alone application which will be 
			put into ROM, or for the special case of building the eCos GDB stubs 
			themselves."
	}

	cdl_component CYGBLD_GLOBAL_OPTIONS {
		display		"Global build options"
		flavor		none
		no_define
		description	"
			Global build options including control over 
			compiler flags, linker flags and choice of toolchain."

		parent	CYGPKG_NONE

		cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
			display		"Global command prefix"
			flavor		data
			no_define
			default_value	{ "arm-eabi" }
			description	"
				This option specifies the command prefix used when 
				invoking the build tools."
		}

		cdl_option CYGBLD_GLOBAL_CFLAGS {
			display		"Global compiler flags"
			flavor		data
			no_define
			default_value	{ CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
				"-mcpu=arm9 -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions " }
			description	"
				This option controls the global compiler flags which are used to 
				compile all packages by default. Individual packages may define 
				options which override these global flags."
		}

		cdl_option CYGBLD_GLOBAL_LDFLAGS {
			display		"Global linker flags"
			flavor		data
			no_define
			default_value	{ CYGBLD_ARCH_LDFLAGS . "-mcpu=arm9 --no-target-default-spec -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
			description	"
				This option controls the global linker flags. Individual 
				packages may define options which override these global flags."
		}

		cdl_option CYGBLD_BUILD_GDB_STUBS {
			display		"Build GDB stub ROM image"
			default_value	0
			requires	{ CYG_HAL_STARTUP == "ROM" }
			requires	CYGSEM_HAL_ROM_MONITOR
			requires	CYGBLD_BUILD_COMMON_GDB_STUBS
			requires	CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
			requires	CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
			requires	CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
			requires	!CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
			requires	!CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
			no_define
			description	"
				This option enables the building of the GDB stubs for the 
				board. The common HAL controls takes care of most of the 
				build process, but the final conversion from ELF image to 
				binary data is handled by the platform CDL, allowing 
				relocation of the data if necessary."

			make -priority 320 {
				<PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
				$(OBJCOPY) -O binary $< $@
			}
 		}
	}

	cdl_component CYGPKG_HAL_ARM_ARM9_MINI2440_OPTIONS {
		display		"FriendlyARM MINI2440 build options"
		flavor		none
		no_define
		description	"
			Package specific build options including control over 
			compiler flags used only in building this package, 
			and details of which tests are built."

		cdl_option CYGPKG_HAL_ARM_ARM9_MINI2440_CFLAGS_ADD {
			display		"Additional compiler flags"
			flavor		data
			no_define
			default_value	{ "" }
			description	"
				This option modifies the set of compiler flags for 
				building the ARM9 MINI2440 HAL. These flags are used 
				in addition to the set of global flags."
		}

		cdl_option CYGPKG_HAL_ARM_ARM9_MINI2440_CFLAGS_REMOVE {
			display		"Suppressed compiler flags"
			flavor		data
			no_define
			default_value	{ "" }
			description	"
				This option modifies the set of compiler flags for 
				building the FriendlyARM MINI2440 HAL. These flags are 
				removed from the set of global flags if present."
		}

		cdl_option CYGPKG_HAL_ARM_ARM9_MINI2440_TESTS {
			display		"FriendlyARM MINI2440 tests"
			flavor		data
			no_define
			calculated	{ "" }
			description	"
				This option specifies the set of tests for the FriendlyARM MINI2440 HAL."
		}
	}

	cdl_component CYGHWR_MEMORY_LAYOUT {
		display		"Memory layout"
		flavor		data
		no_define
		calculated { CYG_HAL_STARTUP == "RAM" ? "arm_arm9_mini2440_ram" : \
			     CYG_HAL_STARTUP == "ROM" ? "arm_arm9_mini2440_rom" : \
							"arm_arm9_mini2440_romram" }

		cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
			display		"Memory layout linker script fragment"
			flavor		data
			no_define
			define		-file system.h CYGHWR_MEMORY_LAYOUT_LDI
			calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_mini2440_ram.ldi>" :  \
				     CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_mini2440_rom.ldi>" : \
								"<pkgconf/mlt_arm_arm9_mini2440_romram.ldi>" }
		}

		cdl_option CYGHWR_MEMORY_LAYOUT_H {
			display		"Memory layout header file"
			flavor		data
			no_define
			define		-file system.h CYGHWR_MEMORY_LAYOUT_H
			calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_mini2440_ram.h>" :  \
				     CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_mini2440_rom.h>" : \
								"<pkgconf/mlt_arm_arm9_mini2440_romram.h>" }
		}
	}

	cdl_option CYGSEM_HAL_ROM_MONITOR {
		display		"Behave as a ROM monitor"
		flavor		bool
		default_value	0
		parent		CYGPKG_HAL_ROM_MONITOR
		requires	{ (CYG_HAL_STARTUP == "ROM") || (CYG_HAL_STARTUP == "ROMRAM") }
		description	"
			Enable this option if this program is to be used as a ROM monitor, 
			i.e. applications will be loaded into RAM on the board, and this 
			ROM monitor may process exceptions or interrupts generated from the 
			application. This enables features such as utilizing a separate 
			interrupt stack when exceptions are generated."
	}

	cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
		display		"Work with a ROM monitor"
		flavor		booldata
		legal_values	{ "GDB_stubs" }
		default_value	{ CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
		parent		CYGPKG_HAL_ROM_MONITOR
		requires	{ CYG_HAL_STARTUP == "RAM" }
		description	"
			Support can be enabled for different varieties of ROM monitor.
			This support changes various eCos semantics such as the encoding 
			of diagnostic output, or the overriding of hardware interrupt 
			vectors.
			\"GDB_stubs\" provides support when GDB stubs are included in 
			the ROM monitor or boot ROM."
	}

	cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
		display		"Redboot HAL options"
		flavor		none
		no_define
		parent		CYGPKG_REDBOOT
		active_if	CYGPKG_REDBOOT
		description	"
			This option lists the target's requirements for a valid Redboot 
			configuration."

		# The backup image is not needed, since ROMRAM is the normal
		# RedBoot startup type.
		requires	{ !CYGPKG_REDBOOT_FLASH || CYGOPT_REDBOOT_FIS_REDBOOT_BACKUP == 0 }

		# RedBoot details
		requires	{ CYGPKG_REDBOOT_ARM_LINUX_EXEC }
		requires	{ CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0x00008000 }
		define_proc {
			puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS	0x00001f00"
		}

		cdl_option CYGBLD_BUILD_REDBOOT_BIN {
			display		"Build Redboot ROM binary image"
			active_if	CYGBLD_BUILD_REDBOOT
			default_value	1
			no_define
			description	"
				This option enables the conversion of the Redboot ELF 
				image to a binary image suitable for ROM programming."

			make -priority 325 {
				<PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
				$(OBJCOPY) --strip-debug $< $(@:.bin=.img)
				$(OBJCOPY) -O srec $< $(@:.bin=.srec)
				$(OBJCOPY) -O binary $< $@
			}
		}
	}

	cdl_component CYGSEM_MINI2440_LCD_SUPPORT {
		display        "Support LCD"
		flavor         bool
		default_value  1
		compile        lcd_support.c
		description    "
			Enabling this option will enable the use the LCD as a 
			simple framebuffer, suitable for use with a windowing
			package."

		cdl_option  CYGOPT_MINI2440_LCD_SHOW_LOGO {
			display       "show logo"
			flavor         bool
			default_value  0
			description   "
				Use this option enables the logo is showed
				on the LCD screen."
		}
	}
}

