# ====================================================================
#
#      mini2440_eth_driver.cdl
#
#      Ethernet driver - platform dependent support for FriendlyARM
#                         MINI2440 of development boards
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):	T.C. Chiu <TCChiu@sq.com.tw>
# Contributors:	T.C. Chiu <TCChiu@sq.com.tw>
# Date:		2009-12-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_MINI2440 {
	display		"Ethernet driver for FriendlyARM MINI2440 boards"

	parent		CYGPKG_IO_ETH_DRIVERS
	active_if	CYGPKG_IO_ETH_DRIVERS
	active_if	CYGPKG_HAL_ARM_ARM9_MINI2440

	requires	CYGPKG_DEVS_ETH_DAVICOM_DM9000

	include_dir	cyg/io

	description	"Ethernet driver for FriendlyARM MINI2440 based development boards."

	# FIXME: This really belongs in the DM9000 package
	cdl_interface CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED {
		display		"Davicom DM9000 ethernet driver required"
	}

	define_proc {
		puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
		puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_DAVICOM_DM9000_INL	<cyg/io/devs_eth_arm_mini2440.inl>"
		puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_DAVICOM_DM9000_CFG	<pkgconf/devs_eth_arm_mini2440.h>"
		puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
	}

	cdl_component CYGPKG_DEVS_ETH_ARM_MINI2440_ETH0 {
		display		"FriendlyARM MINI2440 ethernet port driver"
		flavor		bool
		default_value	1
		description	"This option includes the ethernet device driver for 
			the FriendlyARM MINI2440 port."

		implements	CYGHWR_NET_DRIVERS
		implements	CYGHWR_NET_DRIVER_ETH0
		implements	CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED

		cdl_option CYGDAT_DEVS_ETH_ARM_MINI2440_ETH0_NAME {
			display		"Device name for the ETH0 ethernet driver"
			flavor		data
			default_value	{ "\"eth0\"" }
			description	"This option sets the name of the ethernet device."
		}

		cdl_component CYGSEM_DEVS_ETH_ARM_MINI2440_ETH0_SET_ESA {
			display		"RedBoot manages ESA for eth0"
			flavor		bool
			default_value	0
			description	"Enabling this option will allow the ethernet
				station address to be forced to the value set by the
				configuration.  This may be required if the hardware does
				not include a serial EEPROM for the ESA."
            
			cdl_option CYGDAT_DEVS_ETH_ARM_MINI2440_ETH0_ESA {
				display		"The ethernet station address"
				flavor		data
				default_value	{ "{ 0x08, 0x88, 0x12, 0x34, 0x56, 0x78 }" }
				description	"The ethernet station address"
			}
		}
	}
}


